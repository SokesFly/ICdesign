module                          regsfile #(
    parameter                   REG_WIDTH = 32
    )(
    );

endmodule
