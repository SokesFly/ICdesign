
module              spi_loop_tb();

parameter           DLY     = 1 ;
parameter           DATA_LEN= 32;



endmodule
