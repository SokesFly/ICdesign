module              axi2ahb_tb();




endmodule
