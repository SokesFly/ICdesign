
module reset(
input wire clk_i    ,
input wire async_i  ,
output wire synced_o
); 


endmodule
