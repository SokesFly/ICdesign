/***************************************************************************************
* Function: 
* Author: SK 
* Company: Ltd.JRLC.SK
* Right : 
* Tel : 
* Last modified: 2022-03-25 05:35
* None: 
* Filename: read_ctrl.v
* Resverd: 
* Description: 
**************************************************************************************/

module read_ctrl    (

)()
