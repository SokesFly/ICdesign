/***************************************************************************************
* Function: 
* Author: SK 
* Company: Ltd.JRLC.SK
* Right : 
* Tel : 
* Last modified:	2022-03-24 08:53
* None: 
* Filename:		reset_syncer_tb.v
* Resverd: 
* Description: 
**************************************************************************************/

module reset_syncer_tb;


/********************************************************************************
*Declare delay for simulation.
********************************************************************************/
parameter       DLY     = 1  ;
parameter       CLK_PER = 20 ;


/********************************************************************************
*Decalre clocks
********************************************************************************/
reg             clk_i        ;
reg             rst_n_sync_i ;
reg             rst_n_synced_o ;


/********************************************************************************
*dump
********************************************************************************/
initial begin
    $fsdbDumpfile("tb.fsdb");
    $fsdbDumpvars(0, "reset_syncer_tb");
end


/********************************************************************************
*generate clocks
********************************************************************************/
initial begin
    clk_i   = 1'b0 ;
    forever begin
        #(CLK_PER/2) clk_i  = 1'b0 ;
        #(CLK_PER/2) clk_i  = 1'b1 ;
    end
end


/********************************************************************************
*generate reset
********************************************************************************/
initial begin
    #(CLK_PER*10)
    rst_n_sync_i    = 1'b0 ;
    #(CLK_PER * 7)
    #(CLK_PER % 3)
    rst_n_sync_i    = 1'b1 ;
end


/********************************************************************************
*end the simulation
********************************************************************************/
initial begin
    #(CLK_PER*100)
    $finish ;
end


/********************************************************************************
*Dut
********************************************************************************/
reset_syncer        #(
    .DLY        (DLY    )
    )reset_syncer_tb(
    .clk_i          (clk_i          ),
    .rst_n_sync_i   (rst_n_sync_i   ),
    .rst_n_synced_o (rst_n_syned_o  )
    );

endmodule

