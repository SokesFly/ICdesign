module mux(
input  wire         ain, // input a
input  wire         bin, //input b
output wire         cout
);

endmodule 
