module                  regsfile #()();

endmodule
