
module              spi_loop_tb();

parameter           DLY     = 1 ;



endmodule
